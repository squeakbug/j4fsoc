class systolic_checker_base;

    //

endclass
