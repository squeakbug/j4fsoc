package wb_pkg;

    `include "wb_packet_base.sv"
    `include "wb_cfg_base.sv"
    `include "wb_checker_base.sv"
    `include "wb_master_gen_base.sv"
    `include "wb_monitor_base.sv"
    `include "wb_master_driver_base.sv"
    `include "wb_master_agent_base.sv"
    `include "wb_env_base.sv"

endpackage
