package systolic_pkg;

    import wb_pkg::*;

    `include "systolic_cfg_base.sv"
    `include "systolic_wb_gen.sv"
    `include "systolic_wb_driver.sv"
    `include "systolic_checker_base.sv"
    `include "systolic_env_base.sv"
    `include "systolic_test_base.sv"

endpackage
