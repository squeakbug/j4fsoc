// https://github.com/nandland/spi-slave
// https://github.com/nandland/spi-master